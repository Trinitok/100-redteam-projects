module main

import cli_arg_parser

fn main() {

	cli_arg_parser.parse_args()
	
}